*Vout and Vin with time for INVX1 is loaded with INVX1

.lib ~/.local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param Lmin = 0.15
.param wp = 1.26
.param wn = 0.42

.param ap = 2*wp*Lmin
.param pp = 2*(wp + 2*Lmin)
.param an = 2*wn*Lmin
.param pn = 2*(wn+ 2*Lmin)

* The voltage sources:
Vdd vdd gnd DC 1.8
Vi in gnd pulse(0 1.8 0p 20p 10p 1n 2n)

Xnot1 in vdd gnd p not1
Xnot2 p vdd gnd out not1

.subckt not1 a vdd vss z
xm01 z a vdd vdd sky130_fd_pr__pfet_01v8 l=0.15 w={wp} as={ap} ad={ap} ps={pp} pd={pp}
xm02 z a vss vss sky130_fd_pr__nfet_01v8 l=0.15 w={wn} as={an} ad={an} ps={pn} pd={pn}
.ends


* Simulation command:
.tran 1ps 10ns
.measure tran tr TRIG v(p) VAL=0.36 RISE=2 TARG v(p) VAL=1.44 RISE=2
.measure tran tf TRIG v(p) VAL=1.44 FALL=2 TARG v(p) VAL=0.36 FALL=2
.measure tran tphl TRIG v(in) VAL=0.9 RISE=2 TARG v(p) VAL=0.9 FALL=2
.measure tran tplh TRIG v(in) VAL=0.9 FALL=2 TARG v(p) VAL=0.9 RISE=2

.control
run
wrdata /mnt/c/Users/anujy/IITB_COURSES/7th_SEMESTER_AUGUST_2025/EE671/Assignment_1/Q1a.txt in p
plot in p
.endc