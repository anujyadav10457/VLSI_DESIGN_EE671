*Vout vs Vin and their direvative for INVX2 is loaded with INVX1

.lib ~/.local/share/pdk/sky130A/libs.tech/ngspice/sky130.lib.spice tt

.param Lmin1 = 0.15
.param wp1 = 1.29
.param wn1 = 0.42
.param Lmin2 = 0.15
.param wp2 = 2*wp1
.param wn2 = 2*wn1

.param ap1 = 2*wp1*Lmin1
.param pp1 = 2*(wp1 + 2*Lmin1)
.param an1 = 2*wn1*Lmin1
.param pn1 = 2*(wn1+ 2*Lmin1)

.param ap2 = 2*wp2*Lmin2
.param pp2 = 2*(wp2 + 2*Lmin2)
.param an2 = 2*wn2*Lmin2
.param pn2 = 2*(wn2+ 2*Lmin2)

* The voltage sources:
Vdd vdd gnd DC 1.8

Xnot1 in vdd gnd p not2
Xnot2 p vdd gnd out not1

.subckt not1 a vdd vss z
xm01 z a vdd vdd sky130_fd_pr__pfet_01v8 l={Lmin1} w={wp1} as={ap1} ad={ap1} ps={pp1} pd={pp1}
xm02 z a vss vss sky130_fd_pr__nfet_01v8 l={Lmin1} w={wn1} as={an1} ad={an1} ps={pn1} pd={pn1}
.ends

.subckt not2 a vdd vss z
xm03 z a vdd vdd sky130_fd_pr__pfet_01v8 l={Lmin2} w={wp2} as={ap2} ad={ap2} ps={pp2} pd={pp2}
xm04 z a vss vss sky130_fd_pr__nfet_01v8 l={Lmin2} w={wn2} as={an2} ad={an2} ps={pn2} pd={pn2}
.ends

Vin in gnd 0
* Simulation command:
.dc Vin 0 1.8 0.001

.control
run
wrdata /mnt/c/Users/anujy/IITB_COURSES/7th_SEMESTER_AUGUST_2025/EE671/Assignment_1/Q2b.txt V(p) vs V(in)
plot V(p) vs V(in)
.endc